module TxController (
  
);

endmodule //TransmitController